`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: Joyce Tung
// Create Date:    2/25/22
// Design Name: 
// Module Name:    KYPD_Decoder 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: Adapted from Decoder.v in Diligent's nexys3 verilog example code
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
// 	Code source: https://digilent.com/reference/pmod/pmodkypd/start
//////////////////////////////////////////////////////////////////////////////////

module KYPD_Decoder(
	 clk,
    Row,
    Col,
    DecodeOut
    );


endmodule
